//----------------------------------------------------------------------
// Created with uvmf_gen version 2020.2
//----------------------------------------------------------------------
// pragma uvmf custom header begin
// pragma uvmf custom header end
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//     
// PACKAGE: This file defines all of the files contained in the
//    interface package that needs to be compiled and synthesized
//    for running on Veloce.
//
// CONTAINS:
//    - <ALU_out_typedefs_hdl>
//
//----------------------------------------------------------------------
//----------------------------------------------------------------------
//
package ALU_out_pkg_hdl;
  
  import uvmf_base_pkg_hdl::*;

  // Parameters defined as HDL parameters

  `include "src/ALU_out_typedefs_hdl.svh"
  `include "src/ALU_out_macros.svh"

  // pragma uvmf custom package_item_additional begin
  // pragma uvmf custom package_item_additional end

endpackage

