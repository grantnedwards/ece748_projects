package data_types_pkg;
    import uvm_pkg::*;
    `include "uvm_macros.svh"

endpackage