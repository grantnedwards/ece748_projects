`include "data_defs.v"
module Controller_Pipeline(	clock, reset, IR, bypass_alu_1, bypass_alu_2, bypass_mem_1, bypass_mem_2, complete_data, complete_instr,
				Instr_dout, NZP, psr, IR_Exec,
				enable_fetch, enable_decode, enable_execute, enable_writeback, enable_updatePC, 
				br_taken, mem_state
				);

   input			clock, reset;	
   input			complete_data, complete_instr;
   input [15:0] 		IR, IR_Exec;
   input [2:0] 			psr, NZP;
   input [15:0] 		Instr_dout;
   output			bypass_alu_1, bypass_alu_2, bypass_mem_1, bypass_mem_2;
   output			enable_fetch, enable_decode, enable_execute, enable_writeback, enable_updatePC;
   output [1:0] 		mem_state;
   output			br_taken;
   
   reg [1:0] 			mem_state;
   reg [4:0] 			enables;
   
   reg [4:0] 			prev_enables;
   reg [4:0] 			state, next_state;
   
   reg				bypass_alu_1, bypass_alu_2, bypass_mem_1, bypass_mem_2;
   reg [15:0] 			prev_IR;
   reg				stall_pipe;
   reg [2:0] 			bubble_count;
   wire 			control_instr_dout;
   wire [4:0] 			enables_temp;
   reg				inc_count, reset_count;
   reg				br_taken;
   
   reg [1:0] 			mem_ctrl_Cstate, mem_ctrl_Nstate;
   
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect author = "BobOden"
`pragma protect author_info = "ECE792-036"
`pragma protect encrypt_agent = "RTLC VELOCE", encrypt_agent_info = "1.5"
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
DL6aY6jN1OWP2iibej7s2OMLmC9VCPUH4qhGEMRtijmSP1ExH8APH6COIlmdw6jN
f+i5NcyDKH/9Q4A0TicausSEe+gt58FEawazeF7j6F7PBIM6FH/VXuGVpcGBAis4
m826cmjAdOUexs0+wUZcRbDZEp4PAKJtjUc+OVL+PMg=
`pragma protect key_keyowner = "Mentor Graphics Corporation"
`pragma protect key_keyname =  "MGC-VELOCE-RSA"
`pragma protect key_method = "rsa"
`pragma protect encoding = ( enctype =  "base64")
`pragma protect key_block
IG/6SVuUe2CcXAdcxTfzb4oQJBBxRr+x+7JTopP84bIyRo789JzIsf78VBfdXY+i
lL2u+LK3vU3RFuVFFpCi74z4JdXbC6Agnsi/nLft7EzNYPTbwFLgN2PB38kWDWlD
g5wAZPmLDY6y0jM6b7R6VbxlY3tF0w0r0331CrrZYvc=
`pragma protect data_method =  "aes128-cbc"
`pragma protect encoding = ( enctype =  "base64" )
`pragma protect data_block
3gmQDUCsaJdsRuO2gP7hlOiDBJ4rcSoWTT1HCzH/o7uV9DdYPsW3YW8olvfxHtGZ
bJsiHISL0L9BODgigxVLlzbcuUvWT5qAm86xb15P+E4LaaGs9dIkv4pXOlCspUG6
wyOG8uBXd+3/f37ZGep7ThRO9ylm7c63m5QQ8JKk0JSNGYFDjVqLb849NGqxa1if
u+fA/enZqndXnNzUvjAZjDJBjvNvN+A6ovrGaf1TfpiVrVr9EPrOTm4DWCmkHOMB
OSMzlrxNtLUT6I9S9tQGgnj8IS6VH/f2scz2eCDWY/FEQzM+UstOAwM8+8jQy3+1
msXcG9II2VdhGFZP5bN7M8HnIJgRXlwqfk89qHeGBJX+IofaONsmhvsSg47BZ3ri
MOY+NZa+ZdApI5yOjHIFliTFst1ryTzInU1epq3X2MdiiDfk8a4kCJDPP6KhwaR1
uA7RidSAEU4lk460OM/RYTZSjcCy8YDM1U0WVQmkC3tTY/pN9Yj9APRxF0Db0ecZ
ns5TUlQDtpeXI4iI4q2uZYy4cE6VKMJZ4R0AppK36FojJrBy0fgBiZ/26NrSrkt2
XyfCSbfDOt57+4zHRK8/J3kM4SHAwryjw3vEBYSvK5orjfmYiZYAEaBjo5+efBUG
0RUZrXrsSIoWB1Y5l4/m2VfW9PXKGKf12Vjzv8QUfpatlq/vOkt44HE6icr3Y6+K
PywBoiLGxekNxC3U9o6IDaUyFbTFupIWboultJmucnivIPn6RA0aRreOfSFtaN6E
h4TspU0IchgBPxGcrzxJah1IVFUT3tMzujmA8I2kW3RLUFPQ8SQ7aNQphFVqonFy
xrxQ0dFUwYYMOh9UaN4SvFPeCe0nX14h/71xQ6lrZzpBBwWk7QrJmRisUBi8w4xG
0pwPavt8klu7LwW43pe5gEM7JihFFDt0O2LshYojWgQe0u+XfHmkDZuFYsxMyQDk
Np4rmgKoFCO9AjVJ+JPOgXFhU9g5PeeNDB2zkGN0widi8R/0VgKK56upNlgf0ImR
pDRyL/Go8eeI51zJzobkKxtAlmBHiMYy2qLU87BHnp2GAJ166r19NJG5Ff43Oxl9
iMxMN5cq3NDObZWZzlaT+G8Z5B63sCE72QVWOCh4juZ6JbzY9j8QJLLwV2nUIvnr
LTKeh3rB+IONMWVs4SJPQltO1erC7UvDOyKcwo/+pFo+Ym4HZZg14Dy9sTEOTZMy
SfoF+bxA0fCwoQR027+CSbQkVpDMjTr2m717LsVGMKXZVmGk20SWq5SopxiLNwHd
ijtF0ZFhzXSUH+BSaPR+cQQ9NVUbnyfGne/8Th1tdYY3VsRWXn2fZmPYzasQKCiE
4rB0E0QNJuKsc71ljnenIrIytcV1vFYlHVaYz8fni0hFtbWkWKAEhrzpjvmfw+tg
EFSCaw6njkPLzF6wBF9ovSfFJDehajbRgf/9EdYoLp3BdpJOXmhsg06O2QBWGV1Z
asl42c98p30JLijepW2NwQ0aI/G/92jz2ToaxLmV9u+WDYG2lGMyDgTYpl+ynXes
5M8A4J1cNZFVkAWWezBvXXIEiF3MXnBuDeyBBlOKMd7koxcgJ4N7DYcoNcy3LHnl
OlU6aMBpts0cZnUQR2PzEmYZXHnXrtVlacW1WsUj5szfJCEqPbPxfYgSkFKEybej
V4OrdkEpZeGNEq9BihXzM4g3EsFPaq81ANL9uMcWukgKuAy64ujtK05oPCXkMxza
PRRMn8ZyrbecLVnUV2faFKYBsrAWZOscXCFu41AWYPP31xaSs35jZ61y+DSQtFr/
sYRWJTlvChK7T8uksJsdnceO3OYgYp6raKK8LZRL1QKTeaSLEozG99h1XDiHU4Q+
MMt5LmZM29ypQZ7M2gT3t6ZJOcII8w/DNcuwtldvkFYIVuwb7bhyadY7lgwDzXEt
vwV2tgibfMp54BQorXkgw+TO205VQqOyNKYV+Ucg7bxGRaomP5xwQLWxFb2iD4ck
eHJ3DWz8emQP5aWh1F3IPc4E+XcE44VJC55BSJj5Ndw3e89eIdVFu8W6rqwmI82+
DbwC77bHsurtOdpMIHGziROjrWAvyt6ILVZbGidpsIx+YUehy82OLpQpwXDgazuv
1v3yAqHvKzER2Ru+bxHDx7C9oQNI0QDasuBBZnygEuuNthOKI7i1YijYmBO055bm
05LvuO5F5AEmc2yhbsZ08KsD/KnrZZntv6dF3swPBf14L+MdxMD/TNdG7osCKluC
yhbb0uFFDtx6O44iN9e5CaswDCf+v0EEjWSba6VfVDogdWkB+WylDEQrQ1G/lfF6
QQuWb74aZ9HgedFKz0aC2CuJ+NWhsenDC0bgiXsZg4qwZeH9SGMPQCLwL++/+4ZV
nTtMROufBZjGwg4+YTmWOjdBtks+dDWlAuC8STp31Zo8BpzsQ7Kyp4ruIuialnGn
+FvNDyk4ej2Mt8nwukcJZGqfH396sKPShCb8pZAgHIobGzJeGYqQKI5qbz7+mrdB
41KbYYQ4mhRfN8ALTVeLaWnDmAn4lE9IjWnI11IFMmsRPGw45lOD+HjJfmDLjvVF
R/r7sYLjgfftXjAQLTHobyE+RiDS/3aIj0jq4nqLwBUHJuJ8Qy35O68zyPEyDQ1a
s57ZrO5PiSW01NAXf38YdtHFTsxfN1YU/lhQFq1pKleqSDvsnvkTYYc8EiKqzA1B
v8L+QtEmPNR1UNv7b0RKPUbU4lCuaDKWXg5AyJuPnlxF+BNG136IH2KzduorpKkZ
3Dig42YqaxklKeG7SplYJSUMXjaProP4hivhXeEHNTncVACItcHGqzLb9/NN+SEy
UL03phBDyBnJMD/gjiHo8WtZnJtyh42B3FR3LyWbEzhJBCtQaCjGikOy1+YM0PB7
y9a2Gz1fQigjVwBrFR33ud/qewIZAoxZvTuhb8sW5X+TJTWWrfGB8mSp9rZn5G89
mliWNbZjOtD7iWXbW2LAO24KYVV1ktyhbmaDYaXAjgPfNHM31zxEPX71smYNdkhV
NFUZyHrwxicRtnrU0zVUe2sbCqugJlTBH6T5QsW2rJh6MmuqayWE+wjl2fnWg+wA
nctSOfaGlszLoFAKJ1SV26g0t71aRqnBxVnskEXyRt4wq6+O0PNJfjr8z0f9aYeY
OFxKxqgnvFg4NpkOVb54K98V5Gnv1J0uTwjmc6QJ23wYh3zHyrFzi8ZTVS0h23h1
jfpAuF1jUm2oB7DGwXP5tIPnXoVVbT9xD2mxHg82L9MOiMOhfBf6uwM625V6nbSA
f4T6RJhEftBbjffLPDVvgbUQHp9hPhYTsoRF8fOloS0rlb3JlB8nxtS1tkxQpY34
k/9PHQsglYZPFb2FgboZaRM2bNG2vLOSihIHKl4/XDZUppAk5g+Qio2wrmjAd3+F
yoQSS7OvU1oMMMBFzM6J9a531POliHZa36HytrkbOxWw3yu+FmayTKqVGqRPOxs9
AEv9rSJussreEY5Gz1zrLdfxxPYrX2gPYL6Wz9XtmgWXs4CYIWlR/FpTCkXTHeDL
db8qhfUAUca6kTEwXwb2nOGhJL4Njd0nwAWwrG40y025xTqQTIat//82Jq4TogOm
yfzyW2+RljVvItT0HKm1VdKl1m96rIchoeA7RzwcGndUvf+k9hi0YEq/YHT+gUt3
W8+mVOgRMR8BuJmS9V/pQBydciPjEdLYf3pkrwg7tgwwm5dHi0KBuOyUUq6iSYm9
4ThqAO/1sSui0Vs2xbrbM/hJVMdHjAZKqRkxXk2pY4hbQDh/j/d8/nEpjVJ3RjYq
JKdkz7paYhYjhNbOxj/ufe65Ok18p3WQkN/ajosAieLNBIhZYo8V0MlPjaWBtUbb
6WOwqpdGvjQ3kW802K8vg8ALfXaQKsNdlbk9zDfDc6iMBVuO0F3j6aRgf9K05m/d
hR9ePorrUtAZpcydD9P0G8UKBf5ysiOv60od5d8kQkjiVKa3MVswiW+06u9mfnlw
3wWx9+Cx7UtQCHxHG2AN9kp0OmXEacHHexGNuns7C8ngWTtKpgRBQSs5xiWSNaNm
r99oxE37o1ltEqy03LkSELaE94ONk7HBy8uyOWmMogmd5jo18e8uR3GW8IcmcYF1
3IjK4gYO9nhM0lMOjN29E1V4pByX7eTpADfYRisl6X8jA3v5/lESORlVZPhUBAUn
oUZXAnM+pVwSWkVPLzDpftC3gGf3fsfL/yoUYKxdnu67t94sxbH3zTLmffzNTIBv
u06LyWLeO473Nc3YM2/v6BjYrq4kmmr4iH0kOJEESH8omVmGZGcLzdcwFvLefTr7
xXrBuOwCU5p+Ie1I0ZGKr/TnXpruoDlKyKNMyLLQzTju3cPNmiokX3gN0/5ZoFLk
edgcbSzuI2EUkRn4Y3gSL8QcXa+8rE0tDOXK7U66OwAqO4KA57zidAupiHbe9maf
+NkMaVmiXBXN4fX/XwaFnPfaN1CaI1Z4GsV/lxOi16QYDzSuk3XJABKtoaB4iSwZ
V2DS7JfM8w/OuSsKREPatES8CryXyFT0kXOic47ca30bjk0+i+Ph+whZhEbdQ3L4
ctfYFIPm5gAkkvGapbZPAdl/pLfRPoIyXV74QpVGhGYxXjqSkO6lboC3ySloyFke
dAlc/y7Dw5xmDbjW5ZQ6xubpZqnTVlBGWetNGwJ52iXF+u5CpBR2XRjtCScDvFor
VGEoxnvRiI9mPW3YzKfGT8vudHt2YNaSs0SsRVWuWvH+XyUKQdzUXanYN+QzVFJq
yuY/wKVH1MDZxiSOUaD/Mno23suSuwemKfK7U3Qnxg8UzaC/dZ3fx/ClPzDX4mdv
G7ENFWLFGxZEbDnFotxCnrG9j5w5OHsd47djdNRlv4l6qLeEE/NVKNDJmwwMVKrj
CgR9l7hZqzuBHvVbLj269bXmeng1vvSawMsitLX29oML86UQiWOTL4YsPTIkRy1P
Yxv8WZtFQR0AJ4C8yiW4E5PFokWJAiGc+2eDMriv8Ed4mNeehpFEeLNilQHE7HaW
BIER1kuxkPfIarj5dFfUgvlb1a1Y5NWCmxxdxVOMQsS6MiCQ59/73mHlhNhXCBAC
ikacP8p+B/HhO5x00SztviILVZGnAxgsEF0/3Sce6fuFu/iPuxQTdSNljZDFuNoY
EnUPft8E8Cq6uxhnW6ycPrtyoEhHJDQjZXNnsuzR20xxv+PIljR8bliVckbuBnCH
3tqt6rmZuV6vkts4XFtyPL7KTESy5UrndlouR/k6Krff38SCLlDiOks69jBiWfP7
8y6cIw6tjwpDv8igfRAb1SepbOfgcVVudB2KTTz57UAz/32+ImzN0Tx1TD/phd+0
XFnR2j40roKj2lLD49nY+l9dGEivI37cMTIp7pKdmp7ArVTiOqo3qelnmjBtKnE0
Foj62xArz8z5lIZaN6kaiKGO/bm5w327sM2lmmxTCdAYcZf0ih8ap+1JZ0I2o5+N
vSi0X4u6yuHzdYM0vnksc/FkxDtUDTACJps1H3Y46hoSpU3e5mydD+VNDLw0WIIk
AhjL0K/0l9qypl8XO4j/TEabXAOoEeyPLuZ4W70K9tRwL14bMtRB73/MotVALHw+
OyusWcNWWRjATWTtVakG5VAMtbs/ayYB1STRvysN4o0iqmfSfqSyMooVq971l5pu
L4BoD4F3hVPIPSvuy7pjkcQsTTmzifd3qyy6ApS7vhEmvTal0wXD3TaizFtqAmsH
uo9o17ejUtr0IVPgIQjOdN8H9HfbkuYAtI/dGBCAGpytqTFINSdzQPlZIt9cKjs3
ObSiIyWJ5utJgXVM7v4qivYxP6dxyfNZCBGNaRhkwThJH4G/9nVtp8kf/tXMj8fL
lGICZqE4VKpTSCwIY/q0eBD6Ac+r01ibibUtP1p2gtqhlF7D/p5vSL6KvR7maoxn
p8simpFZyteeE48zKKsvwsCWDZcblZSs2yl0GIVI7Dg+VLWikaDC6R0BYS3U41LB
+XmE6J4D04CdHoZ8cg0rlRtDndZuJX8iVbnBlGkmIlRB/eqTR3DMx/whsYWuawEr
L4kbwNJTnu2JJVAPVv8qrBHwnLXabosz6Fcb1YxSm5tFViJzMYJZDSOUmum3b98X
RH55Ar54oxZvOorLOx/sEkgvKYJmZRMxMYJHqVpMxm+O8mqWJA0YLwI4kfJmWamx
/a1wy3kpTbnN+Jzt9hcFFzzn8z73S3ZABsXF2F3itg32VwJre/CbUJ3O1yCmRwKG
jNQ9GXzFxRoTC21N0UJpiOGln84BLc72YFQ0vks4JbS6eQXJSPBatyD2os3/mVBD
PvX7LVfMOX9AuCbxSm8Fw/HWfg4L//zG7GgNq4YevcDT34jkTbyskDvzP04tLwBZ
RwQ2GPg6AVVTxocRMJp6z0HSBUMWTIoaNTYQBilaYGcItfFGLDzrZ6jRLKq+ldGj
hkNTxDGnaZd8JUCxnGeVWVaKjl6Rxw50Iebm2jbWPPgpcfM+2ybMdjbAPKSRbJsS
MnP3ukfNxehmA/JoVyl2W5FTtNsmTFAcmIyUqbAzhPmLbSnteVw+XITLkWIgH/Vg
eO2TkZkZDKAHmujrD90FZcCY/3ZQq6cMnvKYKVulpONmwVEp2v7XHSJO1FDeMjpb
sdEElwpXCjBrh8QngSiAUWekMnxwCIimS6WYXpUYYEUB0pE57asHsRR61AJc8QPY
CJ4psk7TZ+227Y80d3jWJ0bNJmGsCxqmhc7fJ5cxd23O4uU+hxwVFRRDPcI8fNEL
JOGtaSGTm7prooNA9LHqnbNow+UcN8/adND1K5ptmJtsv/g1VDzU5ZiG1T41eb1c
yIY0F6wCVWdqUUhtKA7+swmqRlY9mLobCAdI+D8RxA4UAIzrBb7QdbTX0oTKG+Fh
ps7bG5Z4GmjUk8Be6zWGOGAQZBJtn0AE6OflHXpJQVhnSpp1aYjutSSE33nETGeI
1C2t06HweByQNfIFbqpeklvL9fJr/izTE3oA8zuIgn6EvJKDQoK3j/mvXt+DPOWk
8VixdlKUftDFy8y+E1aviPIlL88Hk3J6TI24segdQ3pl3chvSX/b/jg2i6KeWzEG
ahsK2qgZoFFq8g9el7doBIsNcn0MZn3rAekwuRsC1CMjWLPsn5vIfJOnw6jlFTRR
+smLsR2HJZf1jMCVffH6gwVIG3gDFEyOCplsnZonc9Lge5tyPzg1w/RlYkPDZcLq
sVvG5ZoMj49Vs2/8lvDSNhTsZ0sZG0YLwmHumsNzoN9ap31gs94raLfTvLXjowqo
G9+ZoDeykEFgbvXlp5lmvGOrYXKHbaRVMIC/3nyX/zk/4diMmGv+yZQxrrv18/Uu
b4fWpJIJk3Cx+n6iYdWWVBVhw8xC1w2AVlE7yFdSvSgUPmpR8VHjUteFX63h7jyl
+REMUSVuOaHhYhfMpefVPlAFT/e76jIECMCYpWHK6K6NUVTvylsn5PA6jLXOjBmO
iQbXamtiGpo3P9W/fPLyJJOvC5O64xzBHkeRnKs4Aih6GuRNx7UJ0E/q2d2dIgFX
Tx4eQ97QJsSmTh/XPYmNmZ5gcvv3t6C1HifeAao2sl9nqathI3zE84ECuROER5/x
FHHx+ky0kP4z7N6Ws5jx/FNkzv8dOn3/MJCBiEGmwaEEd8zZwpOG1Kmq8VrlsZGM
MCFi2gAch69acs8OfL5w7Nnly8t0BIipcyLSCYvTHPXfZfDk8z9J7M3DBFoDZEeL
FxU76+/gHl7Obv70VOUztvkFAL3OgfkPHkMBpID5EnV16fAjO2jfGIyaXZYWmi2m
x8xm8VqeGvVrr4Fnw/O6Ot7LH70sGEqETxh5bRMracp90OYYYxIPmtSuZPYj+itu
J7ll2FYHA2d/MFzvBnssqQeuPo7vF5JbNhGba2d3L/pdFlDmkHugX5jJAKD+1f/a
KkgQqk/7Vu3kOFKyolphfhiO/5nqKnvfApmR1/21JWQTthPNnvfFDOkLPMIGqpq7
liUU7Lf45goIv3SARizyWvRlXYdoYJrMdTXsnUw0AFsS3a7+or57DvvL5Q1aQ6n3
VK5qbYVqjYXKoTm5/V9LRHQGSi5rdy+alYUx879rQUql545UdPxI+xZTjc5E3k5I
kphKbACp1ssMtSGfXpvZc8Mfz8L8mYidVUMghK+wQgErPdgzXd1snJ/JPQH1QYWt
8t+4+IAFOGwT9JCk0FxCsImUc2uqBdZ9P03+3Vq4d97VmGew65HlSrks2WrbP1U6
9PQjaNX+0v7y8GVyoqnQdptEM8Id719zqm9baM26brK4VTYAVh175ZZ6DRk+8DgM
abf4QiUeQviOEZpx/gUez0VczUP/lQYOIVgiDec+2h6cvnSth+kzLcTz/e50ZcGy
0R/7m7W+215gd51gU6JjmkNiXyQm5KEPrVUrjiU932Y8+s2n6F09xvJrpBDahS4L
Y+OvEvnvPA1vDqLvEN61ZeeIb1jb6dxNiBd2VrmHG8HVOn9YysQrcRbdfo9eTqAS
A4njJe6kNBjjGyNT/GfEjc/D1zaP1FLKDjqg0hgWmuCRvw36LoLFKsA4LCoPthBc
dvLQ05wcUNyIMS3PoS4vCB2YHw8dhLtKQ/nKzJw+pO7QJjJPD+cGaV1PlXEtWV4+
5uIOIgFpVlliK8jpME0ASMO4v70C+r4mIsQ+LnxWw5gFZCWx6AF5TD6vbKQyCiik
De/0fKPn4vaC8NXH2Ya+xPkQhOGPXt2V2nMz9p37ZvfDMftvP5ni/xWhmr3k8L5+
R46jCH/LI42YjKr7zW++UQIBxTe2JqMVKWPjkh4Xu2ar3xH4LpYVElGPS0pslKt/
ReTBgmBbYGskioF7H3Mf/E4/6aTd3bVq442kZGbjmc1f+zZLppUwlslV5ldsKh3M
rAr9bLurL5NwzRfzJahyD02kZxlLzliTPjuAav05YD1YYy+yrRVR+c9HjDpPOqfp
VxBoieQpUYCKg9UbXLGRVWM1SHsfljfENod3BjZjHWdxdQ+8+a0TgyJezjAYEcrF
XX1chayoP4vEVyZ2KGNhMv3FS0e3ZfDLrZ7IXYKYDxk2/X6C5tk6RgMF30VMqV7g
uegZjbp8DgZ1vRfclyzjxTtJelgbszhLNP2jlFgB9lfWqpQU3+uaxk2yk7xjTst7
QkPJoQ5JW7ycL3AvWlBzq0kQz0R5QrEbeZqYLode3kDtpntH5xEE6RfgAHv53Tvt
FrRw/oymaAm4goYeudqbK/PATXKwCIYEg2rcsgPxnk3Jy+LkEVtr4+g0mh0HLZuN
OaTv1xJZQ2xoGvK/iw4WegItuvTXSJ3941j0zp0Ek6U/tvwtGpPU3ZKT0vplPHM5
CybepbX2t5O80di9MPjuHy2qqKNt2fTxs6a3d6uKjGibYpt3YY9/lfudsbz5N3gW
V9+ilKZB9Oevkm6rKEtVZar86Nxxwfu2OYMLWfcPRG04WAo+Ur4wAl1mGttsp8ka
EIUi/96DJ3vkO58fn5/DHy9ujydNwcUg6YVIUlCOWbQT/l+01upiyBsEJl2eVUmW
EZWgYcf/RK1ZgQ+/VbJDgFYrnFqhJqW5erjv/yd5m8L8jCZTxShQVOXfYvXxCnSG
PL8/BH3p8NzpWfk5iHw7moNBODb3enKv6TkbEKEB/7SNUYqb08rWrSz62hjqFBAs
qkxRmz/AQvGIYN9uwYoG2VHGtWXU2/CHoygNbD1BSK2dLMuu09PYcv52edLeYapT
Y47iqSVFw586jOPAZMHumO0UDnocw73X6fcEGXuGB4Pb73IuTMJGHQz0WJu7x8TJ
Jo4h7LNbN4TBDhhY1+nWWFf0LQ0wLKN3/BgtXfuifP6dMKmEsRRXgiDuZrur27g8
2gnvbfTPYZnMQF1GwfwhDxJdTFWiHiC1FxA9aqeiElAEwGFiryGPzRrSCZegS6pj
erAhabEnKLfFkJZQlKQw26FWHATu3Rfz0XMnN9bwFIUW5iiHqm4OaCzK9ZdHVgjQ
YCUtFle4Hoo3Ms8i511+qihonhG9SXGnTiyZbXcREv4Stdjz1m91HYnOgVKbi82t
BUKI+gWXuvwNc+OyDICiW9EITJiMW1OuHCnAD+pVWf9Ifuou+5tV1Ak9nR6fjO1D
tJQadeRz4wFEH2Pw7N/bPiE1j5Qb2C6/ytyYPUHQ44rDESIyALMiU+/uZa5esBua
L0F6NbAA53yCib7B1LCal6lUyh1Jy9wGoLNPSV8O+65q3iJ/wp9lJ9X8shdmx/Dq
vn+NOm13PCOrY3GzlTHNMemsleM3kCT3QNwNCLS7gWhWE1gwOtBT7PuVkOgCWrlO
MZeTaCtuibE5sj0kbq7spe8N3ibjS3feOYy1DIujYs9qcoiQVDyS2byZA7onSmTq
jzJWthnGmkPHfGILNVKISYJtSIjfSiCSG+LWIAdqEpQrEUgVLsHxBWMoEC4q5mkg
qLuL2vFbciW7yWxUIq3FFBRDeVeF7rJ6EaopdzWryJnKglU3QvwyN3HQZ7uBScgi
LvfPfl+hV54/VEKzUpOVVcCcFrG2v9+Gh8Fph2YV7q32WPlZeDMdG33d6/kISJo6
XlynOrS6QkymrVI9/g++FKHfORoPPkIAqYUsx192smnA7p09ggoEsFB4Mumm/h9z
LmTV1B/f6KyoncsN2EoQjeSqqzathtmchlQ+kAXUXLEZlp0/EAo/AENi+H1jv/lt
YzvOT/ILzgjpXJvQEL5jKNbgMtkn0gCOu/gPGZEV/QaZrEVxI341WFlerA2/AlDU
Ao/0GiU3bPk/L+kbBUkZrz5o+PVL2qZWR0pcJgE3WjPEbjPHhQhsIBMEtHC6Siup
BEmHD4/rfS59DOq3TZV15aaYwgPqpxg7asJoD50kQ9/iVbbsL3KmW7UkhXbU8hKs
36iry1v4U3OIQ+cRgXPs17XQoI39bgoF83WhLFP2OaQLTq98hd8DT/n8TcRwoQBs
snEsGd/z84NzRHvkkAWdpj0oOdnVKOJRlGWPh6UpEwixNpw3DBqmES6FqU4OvhFG
NyoxFksJ8OuKYLWJwH7Qh3hIyFsz8nMpayBa2XSx3EGQeQAw+i/U1tefX2H0skCJ
XdfCbWIx6NpI/b3Fvmg9D3Lmb5WigjSmdE4tdrEItcfGzlLzNyCecvfkR510p9to
1/VQ/giP+g0VSPEeePXRLLVX3WBYFyhOpN0zeTR8FIF8eNtYwSA+AwJH/B6tv+F+
9GYly6kvMbz+4t1gLH4Zq96CNWw0dFdR7Ig+Lr8nFs0a5NE8Hw6UH+x5PQsZpDzj
E610FdflGFdd6ePoCK6S7/k1wm4r2+fhKPCir6JCPC51kzDftjvmBE3GctQiL0gX
sCntBDhvf5J02Jmsm7ayF97QULNqy+1X2EIFyIEZ/W4VRedW9SF40q/ODn0Esn43
83OLX8F639snbQMF8LsvNqNTDEiCMsmqsnNnuGJeLcayGPnLr70GFrn4itkCHyLR
JOU8S8u8rl7zfuWACi5NuIOIyf3WsRhudLM+wJLLpje8PARxBnITtvNw4X+hauXG
wgWbMx5aLBsJwpVpd+skszbqc0WG+g850bYrZk6s4HPUXrTzttWZldORS5Bo/CYR
ulGmKVzyz276qcpKNhyG8yOLvkZIqu7V6aEQ7/32WDoMWyS6ru3CThOR/ukUoaem
6UWuUrRnk5sy5W56dKa6SMdReB820e+zscJyHLuyeUtUKGaKNEka1N1p50RH7Vof
JauEqh2nhwkikokk+ATjMideP9ConIuzFoF5ox4BZeWihoxMGi7d/rXL1vSE3M2c
N8w8RXYLirrxwI8FAaQ+7dnLsA9juX9xM3RbNAis8K5D/1WnHxuFDyThl+LK0o6P
neMajsTPR/z2qwHqA1ZZiHamti40kiiw/Ja4+m4cXWwk81Ied+D4e+JIPp4E6xOg
FGmAS0cTJt+2T2bUAVuY26ljht1ydl/kmeKQfQI3J9pUNrzho9kuwtPHL2tXmnw8
vMnJlCvVq2nLySmU7dbjOSrMVqVIpbKZIrifiK6noBEYRr37uNT+6IfpKYLhrI++
4Irwv23RFsP5k31GbUTkRnoX91ZKMPqsGQsMzYObgdcuIt+jQQmYiHcVDfeFuxOB
7KPfqhlsOETVwy3ioaBzhhiPOnKhnWc4lB3BkXKmPwznVfxwuuUuR704aOzA5EqE
onvh2WHpuRj1tjDyVn6H0gVZYNNfeeHXFinDYwgIQD6wwo1pXfuiQA4mcoWUGc2D
mXCMYNhLSCdTJvD50isr0VIlkwWX/Gn2y22qJQ0VN7UojN2IuHXKTJmZEiuGGEcm
j6eSKNt2uZGDY+ulGWIswPIU397ctKZULySK9OGkHauQvv5sTFYxGBu2ovwo6cNG
q67oo8fwqDDLObG+ITwra6xiY8mBRoi8OVeUumuZkO26gcpiwLFNMyKZ14SQKjV6
7DScrBBvnrRHSa5ZWFkDZ7yz5RLsOZZ8yiM1N4HdHRKY0x5lP9vHEsLI6PXuBBVV
XBT8DuKcTYt8DbBlgrpo9wfLLvRUh0Y/niv7RWpY8tzW2egISddHbW6nFQFLonAa
c0wnOd2FAEMGCY7w4ZXhOdKlnCZTRBczQZhq4/AOXWtri2D5Oxm3jD3xopUC38dp
ZBRn8clzcUTF+oVZzwmtWVrBSjJd+8KO2vcjiFZCkPi0rt6VbwuM0wUlXNmwLJGQ
C5xa0gzQMa6EdQ8us3wgbLYeWhZhyTzdMVegazSo7jKLZeBRwYyO4owWIx7t4mDA
aGh61OWtfCRW3LuD6eYxg6vP+Zlx6d0LOiUKeb7N9pezuiPnwJswDhijx7UVCApX
6RyGY7eccuV7jFAA4pmLcGCbIlYG+s++EU36KnXTRfQ5X5i2NpqDH4gpk0R2fLM2
BCsPCnfctgE5t/2k2tZOrncYj71o+Xq5h/epjqEXpBC5puIunh+ozG2Cg3/8Wh5J
3MfmeKR6ffNZ26gqoJHXfe/ZflbZSlsK/VaHxFYcY40Y8Qw//NiOHrcP+3K7rzKS
QgFeb0Smd6LzATj6Hi5TomimO0K8VXArGNh661Jbsl1Rx37R891hZpj/lHwDZNuo
IrFHmR6FkgP+QosFVvU8M9NFwzjZ8lz+bzRg35/HJcmjC6WSsje4XbQAYMrtSU3I
ZEn5WRBPN8h8D+PMQM1SxHk+5YdtngBv6duQd7xJYfzNTTzu/OMJJM5JkadJEvJM
FreK2Ks5QopuOIY4+xLbEbiV7/+NqXUl74GjKT60Cef5vUhxzG42MrQDtmtQc77D
PFNcnqiHiOCLdUMgf6XRjOuSCeOvWhCPAKYVNjgt5HoJtOxe2/eDgUZABVc4jFf3
Zc5xozb5VX3SJk62MDh9GM4ou/sFmpnk8sdRNMGpQxmRoUaYubqGO86pQpjXU1Aj
knlKi2KxEpXuXqTDH+Kx/umfEyrYtmEO/sgQw1mFVZNIxo9FK76Vj6uPpEC/nH+l
4nUjPkIkvX147nmTzi/UP5g6xnTWAYf4JKHscOVmH8ii/nnUfiWxnNkqmTZ79U+H
BmcRf4LGlngr/zEOoq9oIzBQhxEAaIQzxEJZFIXq3iES4Q2GX6B3ce5nHw65HyB6
pzuwGgukNDJiQPi9vZXhMQh+V6dgUaPRoDchp33CrTGqsgvLm9PdcYeXs4hptgw1
PL6N5D7wlsPbhehWC85GN4+vJv5vaD5obKgjg7yxXfHiZb1lnr+5nwiqHHG6ySmC
rjUe+GuvvsMZQjjvSIl+Ik2Wecwc14N3Gy4NO5M8AcD3rw2y5L10PqcRCwN4NpTa
FAn8dove48gshuUwKGO/Wcm6cWTgUkbBxBmopaxSL1l8o2FZSAMWD+IVrLRhgi95
xweXkHUNYmXlU13uziqAUZ6oyoba0cqjZ6NISQhtJtQwfWwTS1t1fP3uIpe9Wnha
HZWSilr3FvKGHK33J2nKG98MSCdWpyiF8uPE1aCLa7hnGkCVYgldFa7FwS0Fzplz
RQW9GeQfPHYgE4jhGmXt1W4yY37CT6smbi+W75q5L+2omW8Wk+Jp4TubGmdceoqI
GABVIAX9LrdoSk5RjSzKBAuaXyEzqKNXbV2YXUTw1wJ9aK38fXWztKpCfvz/3wmt
QbfHKsvq3Q8ALZEn2I5jhFBDYYhRkxKVW6v1Im6QtIMgLpyJI1vJk0zzEfnx9Mkt
ifsWB6PzxvSrw3rmY/9qBZzH7mfiABaBHejyEzQ9TUOUiPOLawXtoAqLEZsG1zwW
qfJSHScVB1azF/aVEFtqZxcKc/SXgZOvnBH+GdlY+I44A/iOA0tzLD93Oazd66MW
Hg2Z++GDwquLjImRwmr3lEDUE5JBuF5SNE88nC0ZhHhKoKWBRaNiow5W8TFlAQCx
fSnBOVDJHlXJtq6YgTqmGJlQb9g9GOAlesBXdNtdT7Gklqz4p22+pkVckUsGzu4J
z5OB0A1ogb4Klmu4SEqhvkYNlVmndHeotrR3bFm+7mteKOUk4qaEkfxaGJphOuqo
Wo8E9P2WDGmjSLbbxJR8x0HlA8/kycunFYtR/MRVTgBqWXn4O2z77dFMik+7++Sj
+j/DAyLR2oT75R7evYunhexh2AJkekA8d6Vrjr70w2vrw3p/fqgPuRALKUpziwpJ
pmnT+so1WsolpMHbouBvAsNil79B6VJO1UEORI9lzUQsS3naTyjF7vM9EKesWBPh
tilYzTRfTWrnnR+GTfp20ZOvGnTblqv0HgZGd4nmIIUK+pgrXSWeq7BzbzXLw00T
FZXT5rjg5zAHb9fbGmsrXF8qdXvjAesKcnXEJrJpQkBLo1t256gG4XIvEpbjdROk
l1XmLFAHDUpS89D4wtGIxdDVSRJWTn8LYl3YR7VnyOjTjoxcIbOXsxMvqDirxdAg
giApu2whGzxK0qxf9eg50RpYumDB1PpdzsXvz4JC+reHICVKI+Vmuu7y2bkSGNSw
seE/nUIQAHuVrbuXAisiO62dFyjJWA9pCQju34DmF3f8AOWgGfUnZbY/GrkBxIzc
mlJddoYJcNdt6L18hyJI9m4mPabdT9Vp+ym5r0VGViY1REzHeahkLei/OC1NvwxQ
o7OrWi6tLD5/9GiH9NntmGiY6u4GgyUjcnXMlzzNUYJWIulkOy9tx+D8+3sSeoth
X6L4ewemfzspBsw+qDuEi9PJ902te8MIeUJamm0ySS8gqXjjyo6H/23LCe0BTEfn
JMk3P3MPvXwzrB6V4KnMOU2R1FoxkLl9/iiKMP3aFPmDHyzO4eEfhyGUxnNmYPcK
4yP8VSPSODc9O5HSk+hNlc7AHWTwuExYsPCr/8hVbKMgYPL/gNgAzs3AtEFEsSIW
A4qdmybsT37HUXGZa5C5IeqDRMSRUeaE+JHgRmMo4yFRRiqg0TKyOaCTtdOy5Xrn
p4XaewLJmRFi2Jbzg8Hixz9gVa9Cj6fWw6KolbGdCd3p+9urQ2j5W0VFDrhHyBS+
Ircn5ny9MPFjPt39E5k35oDF0+Y3kGdkS+GjoaNtWYYHCdfDOvkAvBo7gR93Gp5y
CeU40gJPBOgRDYuU7scAnQlValzA8uTbJNzRnqmIbb45T65SBg+gU9V1XXwrXZiQ
oW2BR/A269K6o8CLV8pJQEtbpUTKIuBDu/pAQ1cVOwOFAU0JQ+HXPEXlZHoTWv/s
69O+djbgTfzfJR4lzbHflqZ8WK1wZQS8i5nlChMTQLjMvI6XEF26Dt+hOswqDKWu
zBpxKjerBIU6Btc/71Z4weg2S4fvTfqy7eu6ht/mx/zdrD6p2m/I8I0RCI3FlN1I
4fITPwlRnFzBUgpGXrxO67Go5+v3POVt+SvGdAS6UImp0KtsEJUrh6DwxjSTXF6H
quzs442mIOPDe6XBezC74omOYeQVBXS/q8WN2Y4jDcDOPDJfvXkWB/JSlaYfBrO9
mahUQNoVfesCjsXAjeJKlC862XriJG8moZ5mGh2kDIvwzj1z9zQoNzSyL5/KVQU3
vBY8upDKFE7OBu8WxXnJA/xJJ1yc83Q2RTrGSZkL9OzQnynmmsWQcQvzhsUTeEqU
ynPC22nBAMdeUGflx4Bv3HwYQwM4iTJ9tQLewr7kc76XvcYdyzW1zBtZ20+DdJTF
+uY06VGL30DmX9YxioRJ0pcwWRpH682cMQndjUEAVludg106Zf1DZQM9jUW+aPrD
Ny+H5uFdlevDFsDBHhTExwALj++wFM5GuBn4WTSmnO1HAcbtthTbaaeai8i7DlGP
2EK4vw16QAUCe6tvfeipWW+wK1kYTc00W9CQUWiUAb3JIQnm8Bp29msNMinPYKCR
U9Yf0/wTWGcSWA2JG/hP0GPpG2F7W+YwU3DIqGsGv+6DAuGu3VbsshVe0fddx139
IJ2qXS73BHlzRtw6m7Vc2SN+HywnGvOrnIlIJM8eCMrGeTdtc9vv1IR7cRoH4N+F
KSDQu24Jizz1YYhZckPjFYdPPDUMY85vqv1KROYhmsBmX/T78qxFfvh9xmSdrcwo
NDovDkSd3ZIRLkR1qa+5nTp4yjxQXbXtwvOkU/Z7r50xQRa8Mln55i20U1xmLFN8
F7Lg1+syi+rZ3Sbz7BrIM7W3u+/SN0NdvVOCTENGAvOMkc6KHO80TDRWx0c1tRXl
U1T5CVUXnaE/jrnqpZ0RUC/ZQnLuayf4goETzTbFsfgcgGdhzNPEqMMdu+9Y1VL2
JGdepQlLVkY08Vo6jJ143UHcLTI3yO9oD9j5I+GsQyHJ+nxruQ5jriG3qtOAqKEL
xdoeZcc/2yvER+JIZ2OuRDUwCdJgl0prKRQkKRe8fzhTns6JFg9zPCNiukfMgla5
Tr+YIHB1dXULtKajqXjC+peBZ46L7jugWbixYayebVQFOW8iu1IgJ3QAF1l1CCbo
hJMszv8a/jU7jKJxZUE8L76PL7Zp8tBGSTCJeToWNcdyjCz280W8VhqcSGi0HiiI
b9UaKjilsSM8Dg7mB7jiwSbkax8u1kasV1k5ckShhUA/B8ofA2fkbWkPQuPkxzgG
aexCnlPjldT5BYV4kBJmy+olfa3il0vr7NoZ1OIjiULPMd8kiy9+IM2q6W559x5D
BO4ByBTadAPUGoH5fOLHsFxg6HMUgb3MlZEbHN3beduwg6ztcctVZb9c8CpVSJ+i
mp7XHxpuU/CC8GkqfZSnEac9iNlihPysrCUxzzNSiDoaefNjN1L8vIR9Cy1U8SXg
ZeEfko6eKBMGRP1ytWMkjyzaWFXLLnZRX+qz6I3aEkRSltEk0e7VX5gXdou7Lq+x
GsCQE0kaXehu72+EOea3jZV01Bm8O6B6mLH7Yz7iD76KwYVkJ/fkSFq3egwfo5yI
94wf192fpVPHiuSSvENEW4BBVNoF+LLgb4GbC13+K8kPDZPmPp0pKmed8F8tB6tT
grMdonr4RZBdGBRuMQv9RoqsVrAup0kixgbfJ/XKDWd0mFV3U/UHWKzMqMrj0HOS
exw6NAku5u4kG8xUtg6cpE+xUbG9Inb9FmQxyoTc508BukRhklu9e0IRK71Yvj1J
ZPG8XUZ+uzP3rEz/ymy/McSByMOXSEt9+ZEjzlj09hH+FahJiRfhwC300pQ2p9z2
j38eIpLg/W4/XEciq3/b6gx+CIIdsKciyCT18Lo9uc72LzzBWzNafcvRYK1BXMqd
PVMr7Fb+3e6Bc5aZZof1bFjAbJrmsS+S0y+xHjibiYS5Kz80GSAb5LtwkKDie+Cd
UtE9RVDdwUWOG5YVBOFF01NYw9hda8Gvoab8Tui6IxaEKep469JFykiK056uwuD2
1XJ6Jcwk37lZ2/joR9Aig1G5gLj+bdfyiegfvK0CdJYDVLRtc5afw/94wxw6wTSC
FlI0baL31JDhK1ymZeN56pBERFxPP5DL23dGUIFs8paEqZiKwmiymiLCHOfllFa4
NWQ4RGZBozJPqUIDX9kg3z8oz67T9alfCIDOmejx8t2cR7kHSNMxvgBpmMH6SaiS
KugIfk3wYufTPXNW4qWFQg9E+QlxBsiFca4MFjOqjR9F3uoeSWfTujUw5Mm6jnLp
udp5C/eBpHU5wz11THRvtezFUgqVV7YYWW0NEIXfzKQMK3tvKc1HHCTr5IWxLwoZ
fIteSNsLPYQHl6GcU94XGQb+fhnYJVM+aVkiuw0uQsOgxXp53QT6GRS5i84uPVqJ
8faFTsGbPMkaDeMQ+Znb6rIRsu/WiOmgoGwFviB5/PWrrGxiY371Aq0vCDVzN2An
5Cf2yfAloVqWBL+LlbFRjTsdWpq9aDgm6j72hNAjbwu+9ifpYuKe/Pz/smeBU0Z7
obCgQVCjgz84eTjmxxAsdRXNj0C1cVPi/cyRwYAxikdjiN9rNZaVw74s+TcXN5xK
uJb9WdSC/YUC0V13ZxvTF0fdeChrIVDW1wgQAU9ZZIq0vAD6pKP2iIrhk+3ZM5Mm
G8b+q8fYYify53TPFmfMYlvAajqvYs6Cx03vzIoPrNHDqaHPr4pgkXl2SOO+Sxwc
jC8/zWn1zNLgALnf0+4lORJ7PjdirCNJdktgBNIVh70lxTnhhDZdz7gzbPBjgHjT
B0I/PTjxw4wXC7gvy8Aq8bxSXvHTGOOsKtZTBs7vgv7QYjSG521A4c/pVfwId6kG
1xJWOV4YFW20GmiQ6DPb5c6fENcWLIQxd6cbLhlB3eSfrREkyu+76+d7oWveWXN+
wykXJcygOk/GQQRuFvXrVZJTFYh9tKXCRGKzbrmo14YvMH+V4jz/tDyVFtDP4qKA
xdFD0jx1NQadCXyPLk1fVtbkhhTRuftvrW5DtY4k3bEDPvFUiPfXHxBlgG0D12ge
ByCCNcCaX0eiZO4juULT012gC34xKW1bAk9FeieZttEoiK14yNCaxXaxuZpkouDn
Hsunwrlc+WR03UVFNLCMVWZMYVKzZIzMapYJjOQdm2EfTvongw4cGHWIyXZve+Q4
MVXv8ZRScUX5P++AuWb7BXVvVlM3LqS+6DxW+Wc9fLEL6xLHuB3LV2tPoDSTfi02
zplKjvhUNFBGiCOZ0KhP1XCJlNrd1jHw49D4DVNN16f88hkF5FDnbBmYQl4GAOoc
KSXnZq7TcaDVCxcQYXyZIVGMhpgo9McvbgtYvrQGHxOK7FU6IhFvYoWYalm7co3B
+fY8roqLC0I2QrHF1TpyRJ6GBeyAHsmXOhj11xqnbMHjlUBnE4OmrJMODn2U0GHc
/HV3O4pZTXigiI99WrUN3SzSyzYwc6RFwG5udEELOVNEO72kM+tZNEsCz6ikQ5E5
K1BQe5+vjYE/GbtffWMCVbcZ32UZE73itZ3oGzhrkth3SOsDqJCR6kV4OaCrjHLz
mvYp/Kx27lpHUNFrcbotMVZPZysAJePXnzGPwbNVlx8kJNvpNKHfiZXB4za/awaD
Ikvr0SDw6VbqnXw/NtPS3k8NpSiXwfiTyf3UTBsfNKMdTdZBVsWca8/hIGu1JID/
M6udQvcwDUFKKSIXtljrf/nLqGT16Y/Hq/rDSinTv0pgMHDKrOQkyaJb5waDpNY0
2m4q+8eYQui2CnU9XVzYK/zYcqPrhNj7n2G8HmSST0kPL3QdrIglCUkxjg5u7zNf
/EjvQlWfMp5IfOaEEbDUfovNkBRAZTsn8+7bq31z9yWSVt1KV8skbd9CufYrVRCZ
yiHGQm2sWbLrh533fJg3yDzQ4rWEYQ6GcjaU0zMzPgN/xO4jIvNtTnOwwXlNOkUn
DAOgHPb40oZ9jeWZtkPCk0TtD+bdJU0oCek8jrDy+f5ZOWETXYcFKfYAeRpDUeYX
5S0toE18l9zzsAQzTnJYoQTzOc7ZRm3E0xFxdUN5XVkXo5y/x200Qh3QgPVf1hWq
CY4rYMiA/mcJ2WiYIsoKPJHS5gmlhHxZaiToKro6k2JocKn6r+UemuwXlpK2KxS0
x+X+BH1IMdK8ITLVskV68zgE4HJJEzEnKneMrkSrQD2WRfZBo8oRc+dNkrrYt6dh
IsDcyAbbTZzwfkcd9yFskmnyXEb1wErUW8Vrt0x7s+YQNbxVAyP9hpou3r/83Pxy
yt8+QPqoMY03kQmu/CvciGfZ5nojOY8oSd1cYsL8RyuyebFQldpPCeQbAKyQQs6Z
8FNJObmBBUtA0QzUGiZLzNY7iM8Ca/LbrHxhV/YfB4Ojym0DUvawoi819mk2Q8x4
Rc4JEimPB6nCdtWs2sEmTGkRVl6YWpO/bU2EhO2uqxBApZ3uebJJbCsuaksEEHox
o7gSKYWCL3fknyL25eQ2UtnE7oStwY90SimQOAMAEW6yvIbSotf2jaupuh4ZtA06
cK9qbHmmausIl617Ltd5jgQxqQplp38F1+Hi+yDyXyw767LausVdvhkCAzwjqyzp
CLGdN8KRWGnnSDGv+FMpih6Dtp+EEbIpEaFbwKWekVJsk4O7qVjRdOMcPEOoJGHu
4rm4ilQ91OIsK5HNpZ3oL2EZXL/sLFGYIvpL+WfEE8+Fe9E1hIc3gCuF2K/slUjN
DJDTClTaR4v67vnznQVuEi9dQk9cNRU9BzdV3cKTSit2zS0frFc0XnkzJTRLYGoE
7vV87YPgwY1USHMABeqWha2vJYCJsothVPLPdCivkYUiSPAqyYpEzz9JwXh7X/7O
JNBcEd9SfSOTqo7bGzB9Ku0YnjhmhLnrzKpKyMiRdIJAFso9WUK52r68GaRoHtsA
JszATFVkdbYo2N9KwhT51tgGv1QVwlYVJO9zNtG19XMPV3XQ2nLNxJq7YwTXLQ+5
Qijpd/G1sVeMViKzHcjZVtOhpebu9XjFVJWJy3vixT1AgbiT6/LVG0Nt1HZMT2ty
DK56ZXmj1mprihnc4kF69jCQglahMmxBT5zyGCUo3NWinMIulS8KXN7wBLir4eXr
1n5ro9RIKg0UoZBnTlH0OpFRtP8h5zjS6KgoSDuI4eEZuTKd5NgBgaTXG/lsYKtS
RnPHA00BgJDAElRcL87nqBkITdREBO2AoWgOZx34wr20rb0InLrChEOzVJu8DtSJ
D7pnFJ/PYb6TZ7XVy0Tp3xHh0lO4+Da5JqAVSQ2AsST5CEw6n//DNSGRmRaTieh0
hxA5z5dsry+R+ylod+yU+we7yyCyh16jr1HpQSVmm8/QuN2LUyADzpaKh7HcJp3y
jwcsKR724hKwMCIKBow4GGs7rpSr6CHyj7xrLd2qy/meKLZymtLOfRqJFZaaV0I9
yUwcu3hOCgjrCY8B9j3LZUxOm2HCu+s+gQnqBlPnafbb8mgJMCqv7npCGMjaNTeN
icXyz9U14xTo9z/KckSuQPOtnbgcIsEmA7IL6Nv+gYWcDmojpt+M2BBXlh5QSpi6
hKje+xraTYQP4eivU8KOTi/uxedCykzgrwJtnN+ufrHADqG0wfphYfvA8gABdvYB
81armVDmG6RvlqXIYvixr5Z/On3wqXBxEBfdwZl0260B/8a2ecwh5QNprDt2ytgh
7aKS8/8/jqKRAzVA0GePP73+TvMGgcsMkM0yfCuQTk9qcF5ONcZ2xkt/E2bdz89g
JMY6KF4aR/5hIL0BivrVcR6R8Kxdl2Wm8V5vy1TQGSF4PWus4RCkzhz5HM64k3Sd
PrfA0h5SRjz2slB+MmZMI6jba2Sb8ppX1Fa1vmKoNVjEMivBAvhGmZSkkcb0+cQi
5rJx6WNAYfUPmuXXTurIP45to/1FRPjf5doDJrI40QHkDce7CbMpS1Ry6iabPvvg
okxGFSFUoPXzDVkK8p5gT66Qzz3PDbUXQdbpEclQkivXQnoBEL0O+H42kKIEPjsB
mp0Z37xlzmsh4amMU9MOPciEnwdm+W5V172pOixBb6kw85QzdFoRGZ2CGALiZNkq
v+34bzDjjSkwR42wh20022xC+z6fLvNwH4cAHFB6rv20lOlvuX3LPZzCO21YkawX
gF/Pp/EPdp8wygSc7XEgdnn4IIpgeO+Lq9wq+lckO9/W2+iOX2Yd0neH/c7Q9dxG
rg20gHuxzZ4WMrSr7dTGndI6Q4c3RuG+bpK/sIhkQ81RBQTs59lOsudnfuwqteyI
iDDgBERgWdB02vMw9D2KukLTWUyNgqdGBnFIFTjYjDT0kKnt43g62Q9yQkx+z7ao
X+1Y5LFExAuRK121tVWQgRSPV9OQFkcyGtSOZBIrr4WNXwnYFuP3FwwvKwLJ7VIl
eCF1JR8ZMMANxiR2335w0KFqqP2E0qYkby1P20tIEyRK9V+HPIzgLvhD5d5CwSrm
HHHUbBHgM8PiEsi1S7svNkuRDuOu4x/WagB4fnD0iRYmAnV2PWC82ogOMVkOFntL
XoYBI2rvzWoZ0DbdeOkTigV08H8YyF8+un4resdMTrQMZRk/7fEhd8LAhE/k+xNd
oGAOe10vFpGaB5aAYOmP05v4vDAE7vGyQh9YqJeaZ/fuexjoBqZcFDrV10AAlBJT
+ksjugu5NrmDK/e/2QMsLhfopS988Qog0AClBcnNE2q0ajVnRIoikKS9Y4+62fGU
x0LlQzcgnA2nG3J6HDCmobAVhvTQA5dzxc+uldg97va+Aid9YGPqNYRH+NSdUB0a
wwg3wNurvlDX5hIHoulbqhBGVzqSpXWWNyXebArFTxqhdRUp4ljNdCbAIkvITPbv
rGPrlhvLrwsHbwWnaaxvy3N/x/LRCazpT1kUQvjHC/oabUG9MYqkdwbhLObpgdZK
1Ta7XZO+QX2z+gVom25O2bPKhCVkMWTenvVXDVZQ+xDzOtVhfYZR9Q+CSTIvcIln
jQwVIBZRKFrp5x+7Z6B1TNBx35PldC6XZJYKCmQknETC4RFq5Yn4Gp+cim3EUFqI
Hop4vJJsz2pzc+GHsIWwCOO3OIhEDvATVdFdPXRYJnmJfaGpskHD0F4HM7pvQNtW
VQnY0b/eLMnQo78TqX1woatpj58mlJXzJ2XEqR2MtyxfHE2b2MbAGTKzu6kbd+fc
c15Mft/oNQtHZjpWekt4qYuAsAu5aFBEmvHmwWPjqSdXHvnFDYS3PsffPcJp0Zgo
pTfkXxNvEyrAHmdP63lUZKOPin4INRM/txgneryJMVZ2Y85BgK46c+efsXTsgsRO
hNQ5D/+EaAHcQrjphVrb8rgpshVTu28Zl3jp0IzfTNvYKtDJQzm57Z7RPJKYwinn
hVO5d4y1bvOcwkILfg/O49qF3i4gZgABIbxzXvnvT1Plwmb/zO5yg4qZesn6puVC
O6OFMmyXK7eBbIfKEWJ5HRpvmJILvUO3k//8cqQtJNQyZem6J0ogUkxll9hBVRgb
1pIp9U3elo6n5m5fgKJHHrVJDgEdjcUQiSSnKLgteTtu8QAILnJSQYm8U4iHFcTO
L4yuKUAvP5wWivMoojIUh0I2tGrr/GCkgeDdzk4gXB+iXpUo/UQREFcCK5HadsFm
uVbw/hmHiTQAh3atDGNQAYBfEBvOXJSH0QPNRMiWWY7jV9m3Oqa6fVOmG7PKkNxL
xvDzpZBqfMK2wqnCyUpahGt5wWy1C1yVR37lpnhWdghH82OIUxHRMcUJZpSv0f8N
VibjoOdS+afN8bPw/xNhGeJ5nkq7HGZ7r+wQeSe9WJTpXUDjMaU1+C1cV0pZvM74
E9YvLQBoxYN567R+uwXvmjFs9EeFCvhAw+2wRLNVXpMsLHO8cabn09EHAc+Kb8wF
G14r5G0ZPv58liAmF41fvEJqY3U12r1sRLqxpiaU2e6P7zlXFvufrzBFD7lRYnDQ
jDgSZGVH+N3N0aYOfcA5jlmyYCM9qGwNdKop7pBe8YtLEX/8wvFQ4hVZakSwiMXO
KRy1YaLEis0Trt/c02VDLtQOFcdEwdfaMdvEWJaKzien4CCRk6vsR2RjDRFE/jKL
i6mPrFpAIJCfmuYaNOTdukY8n8Lv6vnnBM+5L5DfrptJ8HtvLorxE4FbneOwcNYf
b6E6CJgmkSlc+xuBBda5jJeBj0bzSpl+/Omrew5O9WxASvKA5yklFgM27OnPPLws
jHuWIeMD4I4FRmubrUIRst2xnwLYd/0SFZspDMgKcVBuAc7N5ryYKzjFMKLUm12c
4EOihp4eZl9RALIcW+svvbh4b2j043n6pDY3aH+eRYFStDNsVCpxeXcD0riGBGIS
X53Hp0WW5hF51PPi+NKHjdjfoGk1PaJcaWiETmwElKd/uxtbtOKj7w7tyssKZjAs
Ik4xUT2h8nznZR0QNrsYY8rat+ZQQbGOTTfXL62NjnwjTaAzWUdyMqDNit32KEqs
U3rBSH+BAT+YKV3dDl5QInTM/lo+y1sjqP+YeZ+xL3jpd1ELp20uYN5eL/byz3sH
mPqOuvyeZEjqUKIIZXVUioCqfg6d+pqkz5Bn0pqdt9qpeA5XfHSPEuFN+rxknyQF
xgMighSZEUgNfY/TbxRWwgyEOu0vdwO7xqOZIrfPCw5g9fVe3vJW1T/TyOPJv80j
ddkiO0KcVfpebloKTKpaHur1gq1tQ8TrEQHbBHHuWgjuAZD4uw0oE+rY/S9aPVXz
eDuOBlJhABGDq89n3VPXqanGEPEaVrXL3wreUJKTHzIlnOAKmjDqmGXeRMZ94DZQ
SCf1JGoDWdpdRo5Ow83UtdL+HKTLL3dFh+S9uFb1wRspEVruak8vJQ815gtnpcIh
Wg9Sc+yCdi3eegCSdAwg3EmGBtfCyveu2TwNrlYWZ21TDa0lyxhMrtzwHKkLDfvP
0JxURZf5NR3A3eRFuKQ/Fbgm3MT1EkpOyRNmtWkoMONSiURC+1EF/e7QP7iKUMTl
/8sWoI5GxDqs7BGaYavK/bRpDDDtUvCPvMYllV4OAL2yPHWQ2hl4vcqqBQkHQ3yK
SLSK3ZlfvlzmsCt6o+qabyG4vlQh8F1nFjh1ZclfxnVAgf398YGV9FsyemoMuLFK
cxwXKGd+7UHKSHtyh9/TGldX0hyZmOlNV72l8jmomDczULu/kk9Jz6yR1esAjOAp
4FLrXqXpE7mbZrpjglIZM5uPtrb18DTnkfkA1Fbs0bEcpS386lS254+fdX3lysLB
XsqlFz8r7uClEEwgO0fEq01Lq4qde3xSMddF4gW/xXEKxJPycswcH427kTGS+94p
ZnqqtKMEDPFfyYc/ZcbKCqHZTfCxY+cSEsie3073DFvQoPz2akoxhpm+UJcqwVh8
dWlPRMH9tkdfA1bP7qQPoxpjd7zlimsu2Nlbu2w6S4nDc0ppSZZdnjKI86h3x5RT
A+f+3bOU1ZkrpiLJr9yBIojSVPfRQYyMbIhs/lvrNRv4Jt+zKSMfR8plN6QyrNds
gX3CeSYUN2kHJEZ78hKjwMagMQ2vR9lqoyRUzBG+RDKlZuhKX1u2z3eTtRahkFyS
80Y2sk8unEJcmg+57LvB8AYlhSNV5PXDWvsJU2clegfKKIvbDmLBGa/vn4Sk+8Za
9eDd/1q/kp67udkRZC77w73CNR/1zazmjwaTj2gEqUouurdxRl9Y1bpY586tDjWK
QKAhbjBVi8JEEzwJr/Cg57fCkc6sagTL/kGmZaQYVvim6Tleg3oU88hY6Ghsnvqq
ndUFeMyoI2qLB2A51yE626v3TjFrPV/c/1uolUVYM/1vF9Abu+MwjJwhxe2uMrSk
RPWQQkB801dZ//NHlUis+n5vbxigiHu5pQeF+v8YNMyAKA7SX6ALPSK77iejwcbX
7is5CiIdXD2vfThL0u+59aOOfpTuxtZjIN2J0mutEcq1dwuUMJAorRiGCndSExtb
4+LldA5+zMo3IJQRuPcQ7rl1yofXwYMSvpZErft6ipK1/+QNsCODw8ghfaQ92bHH
zgSTgj+2W5KKC/ICbeW2wf74pEBeOwW7qo4nZZZQgEugLANjMydgRq30DObeHdi5
1Gf1Z5HWJrL9QjWJfvU/ZA//9JsJlwI7ARtpa6wSXAynnYwd6TeE9Hf++lIrDBbd
1Pc/gkUmiyXOr2mMYfqScaX9f9x90SYhRokVD+3MJguyk01+KaGQAkv+5IgsPPTH
7D5pQ0YSZrLnqinhSXX/DcMk8R0E/IgHI3CW2iRrkqu72sMQhaJ6hvOnbRu8SNFA
ECQ+zgzZJ6DYdeS0vWNphj9HO1dEIn+ZiJ+CQmAiW9lJhkLJ8jXQdeo6/HjabI08
Sj472b7ArM9rcj8pPt+wlnWUupFjEKhnlNF8m7poNbCRINYZMCN2gcdQ3Mgybu50
aqDnGJpdqSF1d/mPE9WBdHYtOgMkJVu69BOT7TQpOLLyDm7pg5cLoxz2IIuRO4Px
XkmkUE9RR+yendKWrMKiDM+APjAhaIb98W1Uvyxr6bCsJ8BZyHzosJpGSQsJEzXu
cBpkFUzU7neX45VdSwev/UxZMxoR1b4Z3SGE6QZLlrloz30IWwPYEGVPJVolWQ0d
g4ZMgKCQcw845WsAWXmpg/cKS9Zrw3CUQfblgZyHb5RmtaJmNtYN1W033K2Q4+5+
L02uW7YjrxPErVThaoF2rkz+6Ggk7vtfDWFEHXj7+uDI/VeSSjvS9u0a2I1Wnt3H
v9yoPD5QaIZKe5Re3h+GNtkiE9TaRMKXRg/7T9Wxmrdum4/7frT4tRgG19XEKZeA
wRyEzimew+H0brj84/y1vfN/T8eVABa4b4z3VsDGB4FkIu398bW+zxW3Z+NAtsZ/
OmFn2zVmkTnHO81fQ4KPwMSd/62r8FGm8z+w4zyl71E2nr2ok9e9QnUHNxeAVWLo
XnS8UwzRLObPdas8J564BEWyThqJuzWtwQN9o2pE+CNmvGjmqAWI1IQ+J8gTLdF8
C8eh1Pxkc9eXcmpOBAUQ6r/tK0rcw8tA0BfLAojtvl5R5cam6R/xb1LKUI4nvX82
TL8Q/Qo8vHPG1otDzrYizWvip/bn8lRaJv0+r3qWnyHc65XhcV7ZLVwvEtpfa7Z/
nqonDFhZLV7eAbTLTMQyL4/KR99XXfoRdjI7dj4KFhyMNZPinBW9ZqaSu1zINsO4
m5mAW8gO1jNm0xr+ctgoV8gqUZY+5tOWij0PO56WVT/6R+jfIEPVNi9mPE/lDKmg
taJmS7xxpudmgbhCDlcz1amctrO+vShrxUSvSdtTEHCjM/A5zMUpDbBBJMawmtUI
QXvyvhn5vuQ9NVuRXE6Nz70582GUxT6tvuHn5pXYnvz33hBrs+RtfQ5HnhtPiJ4b
hQKpkZ6bHIicuSntvhLTF0VhIv3gLTX4ODAByjY7RBrEaP1S1h2oVwYc9BFk3qO1
RHOK1HcoCTrMZ9urGe7QVjtVPR6VH/GxV84GPsZpOWgxwMTAmy9X9VbeT6mKPKj0
0q6eye4Uhr02kViFeCGE4eQUFeBsRgkhWm4XBaVW16VTd3YX/KuACWv5UgeoFst5
F8GTcm3Dsnmz8EAcm1ac9XqZKXXSXLwBvv/YnON3L+L6Ouf+ZoXNZ84mcN8YJNgr
qtb/BY9awIbIqBaedUOQ50lP1BHg39PLWFW9dCJadYtYNWE7ucsQpfIcH9e7dGRg
mirV8RfUdSDgD5a2n8dLfBo8qhobrAs2EEnvfGEHVFmQko191pRcuYLtfco4nL54
oxdJVsTBLLisie326I76OAPV4I0nqXRVxbgbtnwxCs0sGNuk39BxIX4U3na2IaCc
tQUYDAFexSWjEkI6OyQWJzX0BxAHv9CY5cfKMkV3WxYC2haF9Z/2Q00QUGRCxw3+
10cD3Jfkods8HK6lChNvRP6l7PXmJCprZr/ZxTbk/26+Va5Cwu2OtVCOlQv9sQzs
mn6gfNyZckX1f8ohUl/53pZGdniCS+Vtv0Xs9aWQ/p5ITEKt0+zMivKdesvDPmr2
MHbllaZ/XH9swZCoCjzTuinP2aV8JF83pAqRadPEo5eWHklAKGEC9Aot7fV65ihR
LkwTNn/8n5qIpMWdR8y9qdBcGgGHkLQEHADKw9yCP3FzaX/NW8B9vN0aWaHpqE9a
LFK4wWI1vZN+5So47ADqA9mr8sEwYAUvP5b2ElHVpHomAkkFpGMWxiavrhUbD3a4
ZZrjdXr/EGRZHxEgEpfLShgWQEnhJ217JZBVyLVgM9dbLhTUwkCGVrO7wxKgbG8h
YgaSieVAVh4qQPs4q4JcAvtsP89UUkVezuKFIvLec38VA8kvcKszHCRwiQYhRvqa
T85hBMaSdSYxXq7EbgeO3fLD8nqAa4Unowlo7exlJHgpsSrmQTPoAjC9Wkzfm3Wb
NrywIrue3TdHjIbmYGkQ3wONm9eHd3s4cNSgx8JlT4qIc9qT2ZScM0lHk7aEc/KA
no2z4cky4zxI8CY/HvW2UStNOnrsOPkS1fjG4Qiw0hygb57+jvpdnKNwUnmKpAEk
FjEJHHBWEaSJob3pGROa3vLiNPf6vUa9IReviPYVI5S/lx3QaxuuhGylt1+FV4ov
bNynwS7uV7r0uSSo8dOneUO7EQeQMaJgDggD+aTtrp7vut8v4L/0nx3yoymmLlRL
4CMxUzrmaD6jVBbl2zheopfcP41y1L+FNw8/0ttsi9bH0EF6SkuQK1k8nfl/OFvi
Mma601Cag3UCDlbT1n3kwawdW6PdoomsHXL3ZjlnhYh/k+SjwDwBMui7L9Z5k3OP
KssLfFz3AKSQ719NUsESByktQgRSWUFyOgIRPhEYDKq+1ajaN+AugfJtHeI2/BPw
zLixUoi24UUAr1nShFWenC+zmUpGAW3GtkEmK9eekoUOFaEvNz19JsaC6+nLIBBG
g/50pbLrMgktMLM+YF9DkQps9lloH9c3ohMSPCFVow+08Cr7PkrbGQXffXRGX8U5
dYiWolPTZLbovaJZlOkheSqXRt/oayMk252cvB/bPfatiUq2n8MgdN98IYSN8A4P
2j28kSZdACZ0IZMCCxd6kkSo+P9QogDgVzcnGhMsiWSBC5XHPmmIuFkoI7kYJRKi
Tgx2mpnCaKPg4XFHkyV6CycKDBygABe4cmB2PhoU6o4QApje2Op9d9wEZAbdeJUB
i5sNRYgzYWXSxNl/q+GNSy8yUDPtE7Z6gJXJsBAgm4VWU3JqB8KLaFGNwpydpUl4
XAsaj8g8NT1jGC4rpLQ6Lv1Ww3jv9sCLaZ/jeL6re4jN8mCMnsDz0pKzUWV6QdBp
IXS/ZsLEQ6MMcyGMhJjEm/XuTSemGyZNOEamcd7Q+LOC0LuBwINN37bCHjkvpSAG
AdFHVIQJE5jchn1wY7VCWSTHFBvXaxzKpZqxnqCIGTV9wcSKooPXbi4qYH2Gqzbx
LzQ7hc33K8kyV3WYD6/Ve2+oQfl4y8mybv94tcf7T7mWxpRdOL4t24a5B/SP8rLl
e5zQ4Nj4vz164JRAGXErQJb+40+T4uRno34TW8Bke3UqXpwxzLJouzqTAZ7KUyfO
BCA8+F/ZubWkIR2Jn9e3K6qVGU0oXl18TuyDt86EFysEMk3CwdWU1b71QEhpGGfw
GxRcBxZQuh2ncEXpHXufm8EowXWsuXJJNZ3XTfzYJil185uuDavOiGbNgxtlNh2M
KMZPh/gWXLoFUbbuuFGq1+g5J1YV8UjmF0mFw8vYoL8EpmZwliqQDwpK4H7jFGDR
lW21yFBh7PdG7t2oQr1L4M0RTRAEu7xuMX2X453rUYXtM9wkhQGfF+boO+8pvkIG
ooWzxGx5Nzr080lr/emF8bNd7W83xRUqKnPc5oGUmr1WkJM1CBujZcc0a1HNv0Bt
UpstBOtAasGNQSnvJQSbOVdROisguAUXiWYzcMw+HteQPZdqiNjFRjeIneJuJ58b
/ACMsJ9H9JXH6oVGdYgDz59f08kb8c+juNK/XfMgVtkpYLPrC+Irdbz9miZbY/Eq
jcRZNZ2VvlGKj602iXXkXHRSmKnEfE0wOb302xdPjE1KbAR/mZ1O6GTcZvqtFo0Y
vyCCdWoQcnOszgz+nLHb48kQaX8Vfavyzbl4708s+6mxU7/zEna0LnPvir9284Jl
vh/6fc3z2JFjbBntUK8F7BAQFQkGNGFmDOwEqj2qtGyW4x/QxEZx09oFUu2DepiH
02FP5+pru3MdhfA9yAR22XzsaZCUIlwJbU6/YAsfTlwLoGZwYYv1Zz5BCkJJ7gEw
IXmvz6YB53pQaDt8H2YEX+6z+RveGdqbvJcwzEf2g8+n9Mmg8vHOSK0ElAHotdnA
7WEpSz5jgJ2/e6swWJINCQIRUqNSBkAfMmHMhjfkOCjFf9jw5FsoCN4ob6WV6ZXg
vWmT3IFRxqD37YEj/dUbG3yoeVFV7iLM9CPsFo5fHdN14L1kYwksVlFBFiyThmdF
iLd0X5ePcEmhR4KjASWhOQqawULqrFMsf60wg331Wlvfn1AK8bxOeC9Tp7LCDf3Q
hPj1rdverM3n7fqXg2CgXZWGe+lzofa2JUsHpOtf+K7j/itBbyv6CeORGN7x3J59
ZXSwwQuWHDlmgiWjNat20F8Ge1gU8g0ujFqD3bD2flaeqheCf1f0X/9m9AEafyYJ
dmTsKSuSplLWdqmR1cTDCcwKs6o4w62zDssP4bn0wd+n/Wx2lislhpsgGVUborw5
ImptorL0vJ5lsN2SwhcL3dvmqeQSOfzsIXSShbd8D76OQH/tNdePgzZSAwnuAoCP
U+10qVmlgKjrFaZmpQ0anljGkD2l+EeYYtIUSwqJl1g=
`pragma protect end_protected

endmodule
