package decode_test_pkg;
    import uvm_pkg::*;
    import uvmf_base_pkg::*;
    import decode_out_pkg::*;
    import data_types_pkg::*;
    import decode_in_pkg::*;
    `include "uvm_macros.svh"
    `include "src/print_component.svh"
    `include "src/test_top.svh"

endpackage
