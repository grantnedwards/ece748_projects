package decode_test_pkg;
    import uvm_pkg::*;
    import data_types_pkg::*;
    `include "uvm_macros.svh"
    `include "src/test_top.sv"
endpackage